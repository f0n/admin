../../PANOCHE/cdl/wrfsi.d03.cdl