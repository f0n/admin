../../PANOCHE/cdl/wrfsi.cdl