../../PANOCHE/cdl/wrfsi.d02.cdl